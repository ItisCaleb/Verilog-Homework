library verilog;
use verilog.vl_types.all;
entity testRGY is
end testRGY;
