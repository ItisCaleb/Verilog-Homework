library verilog;
use verilog.vl_types.all;
entity test_id is
end test_id;
