library verilog;
use verilog.vl_types.all;
entity testcounter is
end testcounter;
